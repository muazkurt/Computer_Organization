library verilog;
use verilog.vl_types.all;
entity mips_body_testbanch is
end mips_body_testbanch;
