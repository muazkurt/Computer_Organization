`define DELAY 40
module mips_body_testbanch();
	reg	[31:0]	in;
	reg	[4:0]		rs, rt, rd, shift;
	reg	[5:0]		zero, func;
	reg				clock;
	alu32 test(in, clock);
	
	initial
	begin
	assign in		= {zero, rs, rt, rd, shift, func};
	clock = 1'b0;
	
	zero 	= 6'b0;
	rs		= 5'b00001;
	rt		= 5'b00010;
	rd		= 5'b00011;
	shift	= 5'b00010;
	func	= 6'h00;
	#`DELAY;
	clock = ~clock;
	#`DELAY;
	clock = ~clock;
	rs		= 5'b00100;
	rt		= 5'b00101;
	rd		= 5'b00110;
	func	= 6'h02;
	#`DELAY;
	clock = ~clock;
	#`DELAY;
	clock = ~clock;
	rs		= 5'b00111;
	rt		= 5'b01000;
	rd		= 5'b01001;
	func	= 6'h20;
	#`DELAY;
	clock = ~clock;
	#`DELAY;
	clock = ~clock;
	rs		= 5'b01010;
	rt		= 5'b01011;
	rd		= 5'b01100;
	func	= 6'h21;
	#`DELAY;
	clock = ~clock;
	#`DELAY;
	clock = ~clock;
	rs		= 5'b01101;
	rt		= 5'b01110;
	rd		= 5'b01111;
	func	= 6'h24;
	#`DELAY;
	clock = ~clock;
	#`DELAY;
	clock = ~clock;
	rs		= 5'b10000;
	rt		= 5'b10001;
	rd		= 5'b10010;
	func	= 6'h25;
	#`DELAY;
	clock = ~clock;
	#`DELAY;
	clock = ~clock;
	rs		= 5'b10011;
	rt		= 5'b10100;
	rd		= 5'b10101;
	func	= 6'h27;
	#`DELAY;
	clock = ~clock;
	#`DELAY;
	clock = ~clock;
	rs		= 5'b10110;
	rt		= 5'b10111;
	rd		= 5'b11000;
	func	= 6'h2a;
	#`DELAY;
	clock = ~clock;
	#`DELAY;
	clock = ~clock;
	rs		= 5'b11001;
	rt		= 5'b11010;
	rd		= 5'b11011;
	func	= 6'h2b;
	#`DELAY;
	clock = ~clock;
	#`DELAY;
	clock = ~clock;
	rs		= 5'b11100;
	rt		= 5'b11101;
	rd		= 5'b11110;
	func	= 6'h22;
	#`DELAY;
	clock = ~clock;
	#`DELAY;
	clock = ~clock;
	rs		= 5'b11111;
	rt		= 5'b00000;
	rd		= 5'b00001;
	func	= 6'h23;
	#`DELAY;
	clock = ~clock;
	#`DELAY;
	clock = ~clock;
	rs		= 5'b10110;
	rt		= 5'b10111;
	rd		= 5'b00000;
	func	= 6'h2a;
	#`DELAY;
	clock = ~clock;
	#`DELAY;
	clock = ~clock;
	rs		= 5'b11001;
	rt		= 5'b11010;
	func	= 6'h2b;
	#`DELAY;
	clock = ~clock;
	#`DELAY;
	clock = ~clock;
	rs		= 5'b11100;
	rt		= 5'b11101;
	func	= 6'h22;
	#`DELAY;
	clock = ~clock;
	#`DELAY;
	clock = ~clock;
	rs		= 5'b11111;
	rt		= 5'b00000;
	func	= 6'h23;
	
	rs		= 5'b10110;
	rt		= 5'b10111;
	rd		= 5'b11000;
	func	= 6'h16;
	#`DELAY;
	clock = ~clock;
	#`DELAY;
	clock = ~clock;
	rs		= 5'b11001;
	rt		= 5'b11010;
	rd		= 5'b11011;
	func	= 6'h3b;
	#`DELAY;
	clock = ~clock;
	#`DELAY;
	clock = ~clock;
	rs		= 5'b11100;
	rt		= 5'b11101;
	rd		= 5'b11110;
	func	= 6'h12;
	#`DELAY;
	clock = ~clock;
	#`DELAY;
	clock = ~clock;
	rs		= 5'b11111;
	rt		= 5'b00000;
	rd		= 5'b00001;
	func	= 6'h2f;
	end
	initial
		$monitor("clock=%h\t|\trs=%h\t|\tR[rs]=%h\t|\trt=%h\t|\tR[rt]=%h\t|\trd=%h\t|\tR[rd]=%h\t|\tshift=%h\t|\tfunc=%h\t|\taluop=%h\t|\twrite_en=%h\t|\tresult=%h", clock, in[25:21], test.rs, in[20:16], test.rt, in[15:11], test.parse.regs[test.parse.addr3], in[10:6], func, test.alubits, test.write_en, test.result);

endmodule