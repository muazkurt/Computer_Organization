module notxxxii(out, in);
	input [31:0] in;
	output[31:0] out;
	not	o		(out[0], in[0]);
	not	i		(out[1], in[1]);
	not	ii		(out[2], in[2]);
	not	iii	(out[3], in[3]);
	not	iv		(out[4], in[4]);
	not	v		(out[5], in[5]);
	not	vi		(out[6], in[6]);
	not	vii	(out[7], in[7]);
	not	viii	(out[8], in[8]);
	not	ix		(out[9], in[9]);
	not	x		(out[10], in[10]);
	not	xi		(out[11], in[11]);
	not	xii	(out[12], in[12]);
	not	xiii	(out[13], in[13]);
	not	xiv	(out[14], in[14]);
	not	xv		(out[15], in[15]);
	not	xvi	(out[16], in[16]);
	not	xvii	(out[17], in[17]);
	not	xviii	(out[18], in[18]);
	not	xix	(out[19], in[19]);
	not	xx		(out[20], in[20]);
	not	xxi	(out[21], in[21]);
	not	xxii	(out[22], in[22]);
	not	xxiii	(out[23], in[23]);
	not	xxiv	(out[24], in[24]);
	not	xxv	(out[25], in[25]);
	not	xxvi	(out[26], in[26]);
	not	xxvii	(out[27], in[27]);
	not	xxviii(out[28], in[28]);
	not	xxix	(out[29], in[29]);
	not	xxx	(out[30], in[30]);
	not	xxxi	(out[31], in[31]);

endmodule