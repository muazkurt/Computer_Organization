library verilog;
use verilog.vl_types.all;
entity extend_XXXII is
    port(
        \out\           : out    vl_logic_vector(31 downto 0);
        item            : in     vl_logic
    );
end extend_XXXII;
