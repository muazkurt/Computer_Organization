module extend_XXXII	(out, item);
	input	 				item;
	output	[31:0]	out;
	
	buf	o		(out[0], item);
	buf	i		(out[1], 1'b0);
	buf	ii		(out[2], 1'b0);
	buf	iii	(out[3], 1'b0);
	buf	iv		(out[4], 1'b0);
	buf	v		(out[5], 1'b0);
	buf	vi		(out[6], 1'b0);
	buf	vii	(out[7], 1'b0);
	buf	viii	(out[8], 1'b0);
	buf	ix		(out[9], 1'b0);
	buf	x		(out[10], 1'b0);
	buf	xi		(out[11], 1'b0);
	buf	xii	(out[12], 1'b0);
	buf	xiii	(out[13], 1'b0);
	buf	xiv	(out[14], 1'b0);
	buf	xv		(out[15], 1'b0);
	buf	xvi	(out[16], 1'b0);
	buf	xvii	(out[17], 1'b0);
	buf	xviii	(out[18], 1'b0);
	buf	xix	(out[19], 1'b0);
	buf	xx		(out[20], 1'b0);
	buf	xxi	(out[21], 1'b0);
	buf	xxii	(out[22], 1'b0);
	buf	xxiii	(out[23], 1'b0);
	buf	xxiv	(out[24], 1'b0);
	buf	xxv	(out[25], 1'b0);
	buf	xxvi	(out[26], 1'b0);
	buf	xxvii	(out[27], 1'b0);
	buf	xxviii(out[28], 1'b0);
	buf	xxix	(out[29], 1'b0);
	buf	xxx	(out[30], 1'b0);
	buf	xxxi	(out[31], 1'b0);
endmodule