`define DELAY 20
module muxVIII_testbench(); 
reg a, b, c, d, e, f, g, h;
reg [2:0] select;
wire result;

muxIV viiviviviiiiiio (result, a, b, c, d, e, f, g, h, select);

initial begin
	//000 all scenarios
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;

		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;

		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;

		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b000;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b000;
		#`DELAY;

	//001 selected all scenarios.
			a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;

		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;

		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;

		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b001;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b001;
		#`DELAY;
		
	//010 all scenarios
		
			a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;

		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;

		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;

		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b010;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b010;
		#`DELAY;
		
	//011 all scenarios
			a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;

		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;

		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;

		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b011;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b011;
		#`DELAY;
	
	//100 all scenarios
	
			a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;

		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;

		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;

		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b100;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b100;
		#`DELAY;
		
	//101 all scenarios
	
			a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;

		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;

		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;

		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b101;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b101;
		#`DELAY;
	
	//110 all scenarios
			a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;

		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;

		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;

		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b110;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b110;
		#`DELAY;

	//111 all scenarios
	
			a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;

		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;

		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;

		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;

		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b0; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;

		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b0; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b0; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b0; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;

		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b0; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b0; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b0; h = 1'b1; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b0; select = 3'b111;
		#`DELAY;
		a = 1'b1; b = 1'b1; c = 1'b1; d = 1'b1; e = 1'b1; f = 1'b1; g = 1'b1; h = 1'b1; select = 3'b111;
		#`DELAY;
end


initial
begin
$monitor("time = %2d, a =%1b, b=%1b, c=%1b, d=%1b, e =%1b, f=%1b, g=%1b, h=%1b, select=%1b, result=%1b", $time, a, b,c, d, e, f, g, h, select, result);
end
 
endmodule