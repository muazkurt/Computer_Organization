library verilog;
use verilog.vl_types.all;
entity regisers_testbench is
end regisers_testbench;
