`define DELAY 20
module rightShift_testbench(); 
reg				c;
reg	[31:0] a, b;
wire	[31:0] result;

right_shift rs (result, a, b, c);

initial begin
a = 32'b11111111111111110000000000000000; 
b = 32'b00000000000000000000000000000000;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000000001;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000000010;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000000011;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000000100;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000000101;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000000110;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000000111;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000001000;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000001001;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000001010;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000001011;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000001100;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000001101;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000001110;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000001111;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000010000;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000010001;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000010010;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000010011;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000010100;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000010101;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000010110;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000010111;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000011000;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000011001;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000011010;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000011011;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000011100;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000011101;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000011110;
c = 0; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000011111;
c = 0; #`DELAY;

a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000000000;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000000001;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000000010;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000000011;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000000100;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000000101;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000000110;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000000111;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000001000;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000001001;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000001010;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000001011;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000001100;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000001101;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000001110;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000001111;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000010000;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000010001;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000010010;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000010011;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000010100;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000010101;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000010110;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000010111;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000011000;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000011001;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000011010;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000011011;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000011100;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000011101;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000011110;
c = 0; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000011111;
c = 0; #`DELAY;




a = 32'b11111111111111110000000000000000; 
b = 32'b00000000000000000000000000000000;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000000001;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000000010;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000000011;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000000100;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000000101;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000000110;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000000111;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000001000;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000001001;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000001010;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000001011;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000001100;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000001101;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000001110;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000001111;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000010000;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000010001;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000010010;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000010011;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000010100;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000010101;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000010110;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000010111;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000011000;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000011001;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000011010;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000011011;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000011100;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000011101;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000011110;
c = 1; #`DELAY;
a = 32'b11111111111111110000000000000000;
b = 32'b00000000000000000000000000011111;
c = 1; #`DELAY;

a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000000000;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000000001;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000000010;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000000011;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000000100;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000000101;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000000110;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000000111;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000001000;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000001001;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000001010;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000001011;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000001100;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000001101;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000001110;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000001111;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000010000;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000010001;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000010010;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000010011;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000010100;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000010101;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000010110;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000010111;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000011000;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000011001;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000011010;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000011011;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000011100;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000011101;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000011110;
c = 1; #`DELAY;
a = 32'b00000000000000001111111111111111;
b = 32'b00000000000000000000000000011111;
c = 1; #`DELAY;



end
 
initial
begin
$monitor("time = %2d, a =%1b, b=%1b, a/l= %1b, result=%1b", $time, a, b, c, result);
end
 
endmodule